library verilog;
use verilog.vl_types.all;
entity rtc_tb is
end rtc_tb;
